module CNN_Accelerator_Design_tb ();
  
  reg Clk,Rst;

  reg [7:0]In0,In1,In2,In3,In4,In5,In6,In7,In8,In9,In10,In11,In12,In13,In14,In15;
  reg [7:0]W0_0,W0_1,W0_2,W0_3,W0_4,W0_5,W0_6,W0_7,W0_8,W0_9,W0_10,W0_11,W0_12,W0_13,W0_14,W0_15;
  reg [7:0]W1_0,W1_1,W1_2,W1_3,W1_4,W1_5,W1_6,W1_7,W1_8,W1_9,W1_10,W1_11,W1_12,W1_13,W1_14,W1_15;
  reg [7:0]W2_0,W2_1,W2_2,W2_3,W2_4,W2_5,W2_6,W2_7,W2_8,W2_9,W2_10,W2_11,W2_12,W2_13,W2_14,W2_15;
  reg [7:0]W3_0,W3_1,W3_2,W3_3,W3_4,W3_5,W3_6,W3_7,W3_8,W3_9,W3_10,W3_11,W3_12,W3_13,W3_14,W3_15;
  
  wire [15:0]CNN_OUT;


CNN_Accelerator_Design instance_name (
    .Clk(Clk), 
    .Rst(Rst), 
    .In0(In0), 
    .In1(In1), 
    .In2(In2), 
    .In3(In3), 
    .In4(In4), 
    .In5(In5), 
    .In6(In6), 
    .In7(In7), 
    .In8(In8), 
    .In9(In9), 
    .In10(In10), 
    .In11(In11), 
    .In12(In12), 
    .In13(In13), 
    .In14(In14), 
    .In15(In15), 
    .W0_0(W0_0), 
    .W0_1(W0_1), 
    .W0_2(W0_2), 
    .W0_3(W0_3), 
    .W0_4(W0_4), 
    .W0_5(W0_5), 
    .W0_6(W0_6), 
    .W0_7(W0_7), 
    .W0_8(W0_8), 
    .W0_9(W0_9), 
    .W0_10(W0_10), 
    .W0_11(W0_11), 
    .W0_12(W0_12), 
    .W0_13(W0_13), 
    .W0_14(W0_14), 
    .W0_15(W0_15), 
    .W1_0(W1_0), 
    .W1_1(W1_1), 
    .W1_2(W1_2), 
    .W1_3(W1_3), 
    .W1_4(W1_4), 
    .W1_5(W1_5), 
    .W1_6(W1_6), 
    .W1_7(W1_7), 
    .W1_8(W1_8), 
    .W1_9(W1_9), 
    .W1_10(W1_10), 
    .W1_11(W1_11), 
    .W1_12(W1_12), 
    .W1_13(W1_13), 
    .W1_14(W1_14), 
    .W1_15(W1_15), 
    .W2_0(W2_0), 
    .W2_1(W2_1), 
    .W2_2(W2_2), 
    .W2_3(W2_3), 
    .W2_4(W2_4), 
    .W2_5(W2_5), 
    .W2_6(W2_6), 
    .W2_7(W2_7), 
    .W2_8(W2_8), 
    .W2_9(W2_9), 
    .W2_10(W2_10), 
    .W2_11(W2_11), 
    .W2_12(W2_12), 
    .W2_13(W2_13), 
    .W2_14(W2_14), 
    .W2_15(W2_15), 
    .W3_0(W3_0), 
    .W3_1(W3_1), 
    .W3_2(W3_2), 
    .W3_3(W3_3), 
    .W3_4(W3_4), 
    .W3_5(W3_5), 
    .W3_6(W3_6), 
    .W3_7(W3_7), 
    .W3_8(W3_8), 
    .W3_9(W3_9), 
    .W3_10(W3_10), 
    .W3_11(W3_11), 
    .W3_12(W3_12), 
    .W3_13(W3_13), 
    .W3_14(W3_14), 
    .W3_15(W3_15), 
    .CNN_OUT(CNN_OUT)
    );


 initial 
    begin
    Clk = 1;
	  Rst=1'b1;

    In0=8'd1;In1=8'd2;In2=8'd3;In3=8'd4;In4=8'd5;In5=8'd6;In6=8'd7;In7=8'd8;In8=8'd9;In9=8'd10;In10=8'd11;In11=8'd12;In12=8'd13;In13=8'd14;In14=8'd15;In15=8'd16;
    
    
W0_0=8'd1;W0_1=8'd1;W0_2=8'd1;W0_3=8'd1;W0_4=8'd1;W0_5=8'd1;W0_6=8'd1;W0_7=8'd1;W0_8=8'd1;W0_9=8'd1;W0_10=8'd1;W0_11=8'd1;W0_12=8'd1;W0_13=8'd1;W0_14=8'd1;W0_15=8'd1;
W1_0=8'd1;W1_1=8'd1;W1_2=8'd1;W1_3=8'd1;W1_4=8'd1;W1_5=8'd1;W1_6=8'd1;W1_7=8'd1;W1_8=8'd1;W1_9=8'd1;W1_10=8'd1;W1_11=8'd1;W1_12=8'd1;W1_13=8'd1;W1_14=8'd1;W1_15=8'd1;
W2_0=8'd1;W2_1=8'd1;W2_2=8'd1;W2_3=8'd1;W2_4=8'd1;W2_5=8'd1;W2_6=8'd1;W2_7=8'd1;W2_8=8'd1;W2_9=8'd1;W2_10=8'd1;W2_11=8'd1;W2_12=8'd1;W2_13=8'd1;W2_14=8'd1;W2_15=8'd1;
W3_0=8'd1;W3_1=8'd1;W3_2=8'd1;W3_3=8'd1;W3_4=8'd1;W3_5=8'd1;W3_6=8'd1;W3_7=8'd1;W3_8=8'd1;W3_9=8'd1;W3_10=8'd1;W3_11=8'd1;W3_12=8'd1;W3_13=8'd1;W3_14=8'd1;W3_15=8'd1;

    #50
	
    Rst=1'b0;

 end
	always 
	#50 Clk=!Clk;
	
	
endmodule