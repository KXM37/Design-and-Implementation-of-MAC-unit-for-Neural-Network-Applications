module SD_add_6_bit (a,b,c);
  input [5:0]a,b;
  output [5:0]c;
  
  assign c=a+b;
  
endmodule